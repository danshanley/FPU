//-------------------------------------------------
// File: fpu_tb.v
// FPU Test Bench
//-----------------------------------------------------------
`timescale 1 ns/100 ps
module fpu_tb ();
 //---------------------------------------------------------
 // inputs to the DUT are reg type
 reg clock;
 reg [31:0] a, b;
 reg [1:0] op;
 reg [31:0] correct;
 //--------------------------------------------------------
 // outputs from the DUT are wire type
 wire [31:0] out;
 wire [49:0] pro;
 //---------------------------------------------------------
 // instantiate the Device Under Test (DUT)
 // using named instantiation
 fpu U1 (
          .clk(clock),
          .A(a),
          .B(b),
          .opcode(op),
          .outp(out)
        );
 //----------------------------------------------------------
 // create a 10Mhz clock
 always
 #100 clock = ~clock; // every 100 nanoseconds invert
 //-----------------------------------------------------------
 // initial blocks are sequential and start at time 0
 initial
 begin
 $dumpfile("fpu_tb.vcd");
 $dumpvars(0,clock, a, b, op, out);
 clock = 0;
 op = 2'b11;
 a = 32'b00111111001011101000111000101100;
 b = 32'b00111111011100011010111101000110;
 correct = 32'b00111111001001001100101101011010;
 #400 //0.6818568476040797 * 0.9440807186626679 = 0.6437279027111208
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001101101101100000001101;
 b = 32'b00111111010000111110110110010111;
 correct = 32'b00111111000010111111000001000100;
 #400 //0.7142341524887571 * 0.7653440973835888 = 0.5466348927570404
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011100111100111100001100;
 b = 32'b00111110110110101111011000101010;
 correct = 32'b00111110110100001000100011000001;
 #400 //0.952378047779891 * 0.4276593294679506 = 0.407293357313544
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010001001101100110110001;
 b = 32'b00111110011001101111010110010101;
 correct = 32'b00111110001100011001100001101100;
 #400 //0.7689466915660202 * 0.2255462033648783 = 0.17343300687269994
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011011001101110100011000;
 b = 32'b00111111001100110010101010011101;
 correct = 32'b00111111001001011100011000000110;
 #400 //0.9252486420221365 * 0.699868989373403 = 0.6475528320111462
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110001101001101110001111101;
 b = 32'b00111111010100101000111101000010;
 correct = 32'b00111110000101001100001000010100;
 #400 //0.1766223450469715 * 0.8224984579536102 = 0.1452716064412845
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110010111100100000011110011;
 b = 32'b00111110110010101101100100110010;
 correct = 32'b00111101101100000001101111010001;
 #400 //0.2170446355273402 * 0.39618833096639205 = 0.0859905518947858
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000001110000010101101011;
 b = 32'b00111111000110110000001000011011;
 correct = 32'b00111110101000111000001011001000;
 #400 //0.5274263958820093 * 0.605500879813176 = 0.3193571467432491
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101000111010101100000011111;
 b = 32'b00111111011110110101001010110100;
 correct = 32'b00111101000110100111100000111011;
 #400 //0.038414115961869166 * 0.9817306823049222 = 0.03771231627338622
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010111111010101000010000;
 b = 32'b00111101111110111111101100011011;
 correct = 32'b00111101110111000010011100100001;
 #400 //0.87368869918798 * 0.12303754036709458 = 0.10749650859461544
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000010010011101110001000;
 b = 32'b00111111010100101111100100111010;
 correct = 32'b00111110111000100011000011011111;
 #400 //0.5360646261489719 * 0.8241153795308879 = 0.44177910283184346
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011100010110110100100011;
 b = 32'b00111110001110000101001001100100;
 correct = 32'b00111110001011011101010000100101;
 #400 //0.9430715669211067 * 0.1800017965075743 = 0.1697545762810123
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110111001111001000000000111;
 b = 32'b00111111000111111101010101001001;
 correct = 32'b00111110100100001001001101100001;
 #400 //0.45227072117777833 * 0.6243482002106943 = 0.28237441077533865
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011101001000000111001110;
 b = 32'b00111111011010011010110101110110;
 correct = 32'b00111111010111110010111111010010;
 #400 //0.9551056727809147 * 0.9128030817837774 = 0.8718234015435871
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110101000011110000001010001;
 b = 32'b00111111001010100010110100001110;
 correct = 32'b00111110010101110011011011100101;
 #400 //0.3161645108533486 * 0.6647499662977739 = 0.2101703479343157
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001111010010001111011100;
 b = 32'b00111111010100111001010010100001;
 correct = 32'b00111111000111000101001001011110;
 #400 //0.7388284452575336 * 0.826486633568371 = 0.6106318345054524
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110011011000100100010101110;
 b = 32'b00111101111001101011111110110000;
 correct = 32'b00111100110101001111101000111001;
 #400 //0.23074599993297773 * 0.11267030337384198 = 0.025998221814749124
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111100111010111000110001111110;
 b = 32'b00111110111001000001101101001000;
 correct = 32'b00111100010100011110001000111011;
 #400 //0.02875351614985744 * 0.4455206415687205 = 0.012810284962441052
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110101100000010010001100011;
 b = 32'b00111111011010101111001011010110;
 correct = 32'b00111110101000011010100001011000;
 #400 //0.3440276020685057 * 0.9177678574892563 = 0.3157374752675789
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011001001111101001010100;
 b = 32'b00111110011100011010010110110011;
 correct = 32'b00111110010110000010001111011110;
 #400 //0.894444707317307 * 0.2359836482947555 = 0.21107432523067288
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010101111101010100000000;
 b = 32'b00111101010001010111111100110101;
 correct = 32'b00111101001001101000001000101000;
 #400 //0.8430938637777994 * 0.04821701705439563 = 0.040651471208230455
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101011111011100110111011001;
 b = 32'b00111111000010010001011011101001;
 correct = 32'b00111101000001111110100111100000;
 #400 //0.06196388921967744 * 0.5355058425240488 = 0.033182024702650185
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101100010000110100100001000;
 b = 32'b00111101100000111010010110001101;
 correct = 32'b00111011100011000100101111101011;
 #400 //0.06660658086670401 * 0.06428060360842602 = 0.004281511222405173
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001001011001100010100100;
 b = 32'b00111111011001011110000010101101;
 correct = 32'b00111111000101001011001011100000;
 #400 //0.6468603667984485 * 0.8979595245983818 = 0.5808544274518697
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001000010000111011101011;
 b = 32'b00111110001000110110101000011010;
 correct = 32'b00111101110011011001111010000000;
 #400 //0.6291338526917508 * 0.15958443350885543 = 0.10039996948305675
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010110101110001110010011;
 b = 32'b00111111000011110101000010110010;
 correct = 32'b00111110111101010001010000111101;
 #400 //0.8550350040848934 * 0.5598250701005443 = 0.47867003110024464
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110111010100001110010001000;
 b = 32'b00111110101010001001110101110111;
 correct = 32'b00111110000110100011001010111010;
 #400 //0.4572489356197508 * 0.329326364898082 = 0.15058412982116964
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110101110011010010110000101;
 b = 32'b00111101101001100000000001011110;
 correct = 32'b00111100111100001100001100110001;
 #400 //0.36259093395117503 * 0.08105539003453455 = 0.029389949574398645
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110111110011100000110100111;
 b = 32'b00111111011100101001001001110111;
 correct = 32'b00111110111011001010011111110100;
 #400 //0.4878055628913752 * 0.9475473742244943 = 0.462218880249824
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110001000001111010101000001;
 b = 32'b00111101101001011000101110001010;
 correct = 32'b00111100010100000010101110011101;
 #400 //0.1571855647694239 * 0.08083255673531375 = 0.012705711082196793
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110011101101000001000011010;
 b = 32'b00111111011010111111110111111000;
 correct = 32'b00111110011000110011110111111011;
 #400 //0.24073067649007884 * 0.9218439956319454 = 0.2219161286867955
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010100000011101011111100;
 b = 32'b00111111001010101100110100010001;
 correct = 32'b00111111000010101110110111111000;
 #400 //0.8134000216254155 * 0.6671915539520479 = 0.5426936244128903
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010101100001010110111110;
 b = 32'b00111111011000101011110100100101;
 correct = 32'b00111111001111011001110101011110;
 #400 //0.8362692391823181 * 0.8856986209379033 = 0.7406825118765687
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110000111111000011001000;
 b = 32'b00111111011010010110000111100000;
 correct = 32'b00111110101100101010000100010000;
 #400 //0.38269639117588783 * 0.9116497122108362 = 0.34888505487962373
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000011100110100111110111;
 b = 32'b00111110111111000110010001100000;
 correct = 32'b00111110100011000110100000100110;
 #400 //0.5563043966036365 * 0.49295330027417195 = 0.2742320882627945
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110001101000001110110111001;
 b = 32'b00111110001101110010011011000001;
 correct = 32'b00111101000000001101110010000100;
 #400 //0.17589463972975572 * 0.17885877049708754 = 0.03146029899909227
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010000101110100000110001;
 b = 32'b00111101110101111010000010101100;
 correct = 32'b00111101101001000010101101010101;
 #400 //0.7613554481189027 * 0.10528692964533093 = 0.0801607775011843
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010100010010010111001101;
 b = 32'b00111111001100001101001001010101;
 correct = 32'b00111111000100000111010111010011;
 #400 //0.8169830173834385 * 0.6907094173784305 = 0.5642978639449869
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110011010001011001101101010;
 b = 32'b00111101011100100111101101000011;
 correct = 32'b00111100010111000110100110100101;
 #400 //0.227246907690429 * 0.05919958353322008 = 0.013452922294485503
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001001010111000001101110;
 b = 32'b00111111001100000101000101010000;
 correct = 32'b00111110111000111110001110101111;
 #400 //0.6462467745419418 * 0.6887407047053647 = 0.44509645891158595
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110101001010010100101001110;
 b = 32'b00111111010000111001101100110000;
 correct = 32'b00111110011111000110010100101011;
 #400 //0.3225807552268708 * 0.7640867307680019 = 0.24647967466997275
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110100000110101011000011000;
 b = 32'b00111110111100101000010010001111;
 correct = 32'b00111101111110001101011011001000;
 #400 //0.25651621234412303 * 0.4736675881131608 = 0.12150341561296416
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101100110010110000111011001;
 b = 32'b00111111000000011010001110110111;
 correct = 32'b00111101000110110101100011001010;
 #400 //0.07489366028669198 * 0.5064043236401428 = 0.03792647338241687
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001101001110111010110110;
 b = 32'b00111111001110010101111110010110;
 correct = 32'b00111111000000110000010000010001;
 #400 //0.7067674635285706 * 0.7241147883319242 = 0.5117807722528819
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110010100111001000000001;
 b = 32'b00111110110100101010110000000000;
 correct = 32'b00111110001001101001100110001010;
 #400 //0.3954010406466639 * 0.41146850004398894 = 0.1626950731107151
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001011000100011101010110;
 b = 32'b00111111001011011110011110001011;
 correct = 32'b00111110111010100001000000001110;
 #400 //0.6729635070282224 * 0.6793142947093737 = 0.4571537301420235
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010011111101110000101000;
 b = 32'b00111110101011001000001001001001;
 correct = 32'b00111110100011000001000110110100;
 #400 //0.811953095185572 * 0.3369314958073576 = 0.27357257088628856
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001000010011101001110110;
 b = 32'b00111110100000110100100001111000;
 correct = 32'b00111110001001010101110100011100;
 #400 //0.6297982678665204 * 0.2564122650170295 = 0.16148800036745636
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101110001110000111010000111;
 b = 32'b00111111000111000000011011110101;
 correct = 32'b00111101011100101010010010000110;
 #400 //0.0971956764857943 * 0.6094811536371327 = 0.059238933033103444
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110001111101101110110011110;
 b = 32'b00111101110101010011010110111001;
 correct = 32'b00111100100111101111011001110010;
 #400 //0.1863922803343322 * 0.10410637348800289 = 0.019404624351766524
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110111000111110001101011001;
 b = 32'b00111111000100111000010100101111;
 correct = 32'b00111110100000110101001000011011;
 #400 //0.44509389716180725 * 0.5762509961242551 = 0.2564858016083182
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001101001000011001000101;
 b = 32'b00111110110111001111101101101101;
 correct = 32'b00111110100110111101010010101111;
 #400 //0.7051737750374524 * 0.4316057225483233 = 0.3043570366971684
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000010010100001000111011;
 b = 32'b00111110100101000110100111011110;
 correct = 32'b00111110000111110010011000011010;
 #400 //0.5361668345961902 * 0.28987020071273983 = 0.15541878795991204
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011101100111011111101110;
 b = 32'b00111110011101000001101000110110;
 correct = 32'b00111110011010110000001110001011;
 #400 //0.9627674869981642 * 0.23838123973030811 = 0.22950570712265567
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000011100110000000110010;
 b = 32'b00111111001001010110011100101010;
 correct = 32'b00111110101101111111101011000001;
 #400 //0.5561553254542362 * 0.6461054063712333 = 0.35933496255813474
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000000101000110100000101;
 b = 32'b00111110110000110001001111001101;
 correct = 32'b00111110010001101111011100000111;
 #400 //0.5099642641311148 * 0.38101043299277904 = 0.19430170508744
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011111011011111100101101;
 b = 32'b00111110001010001101011110000110;
 correct = 32'b00111110001001110101101100010110;
 #400 //0.9911983319822354 * 0.16488466062084928 = 0.16343340057684277
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110110100010000110010001;
 b = 32'b00111111011110111010010101110111;
 correct = 32'b00111110110101100110101111100110;
 #400 //0.42603732900987756 * 0.9829935648354815 = 0.41879195279640646
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000001000011011100011100;
 b = 32'b00111111010101110101001010110001;
 correct = 32'b00111110110111100110100111111100;
 #400 //0.5164659079166349 * 0.8411055501223388 = 0.4344023415976544
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101101100000111011001100101;
 b = 32'b00111111001011111110111011001001;
 correct = 32'b00111101011100101000101100010000;
 #400 //0.0861633229750094 * 0.6872373200969383 = 0.059214651171992407
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110000110111110110000101;
 b = 32'b00111111010001101111111011010000;
 correct = 32'b00111110100101111111010110101011;
 #400 //0.38181702492680514 * 0.7773256315055727 = 0.2967961600208078
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101100101100001000100011001;
 b = 32'b00111111011101010100110100011100;
 correct = 32'b00111101100011111100101110010000;
 #400 //0.07327479618027288 * 0.9582078364603569 = 0.07021248391497291
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110000111010111110001110001;
 b = 32'b00111111001101111001000011100110;
 correct = 32'b00111101111000011101101000110001;
 #400 //0.1537950231712243 * 0.7170547326825669 = 0.11027944922795142
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010101100111101100110100;
 b = 32'b00111111001111000000010101111000;
 correct = 32'b00111111000111011000011100010000;
 #400 //0.8378174428270628 * 0.7344584702523901 = 0.6153421174095338
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110100010001100110111101100;
 b = 32'b00111111011100011001000100001100;
 correct = 32'b00111110100000010001011101011111;
 #400 //0.2671960667296005 * 0.9436195110408642 = 0.2521314218394277
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110010000110101010011100;
 b = 32'b00111110010101011111111101100101;
 correct = 32'b00111101101001111000100010100101;
 #400 //0.39143836529601805 * 0.2089820663946892 = 0.08180359844572105
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110101100111011001110110;
 b = 32'b00111110000111100111000111100010;
 correct = 32'b00111101100001001011110010000100;
 #400 //0.4188725423171378 * 0.15473129962001742 = 0.06481269284787147
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010110010100101100111101;
 b = 32'b00111111010100000101000010001110;
 correct = 32'b00111111001100001101000110000001;
 #400 //0.84880427345889 * 0.813729144895926 = 0.6906967756257102
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010011101011111111101110;
 b = 32'b00111111001001110000110110001011;
 correct = 32'b00111111000001101110101000100100;
 #400 //0.8076161407333761 * 0.6525503813455552 = 0.5270102206163901
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010111110101001000011000;
 b = 32'b00111111011111010100111000000000;
 correct = 32'b00111111010111001111100000101100;
 #400 //0.8723463816321271 * 0.9894714222539233 = 0.8631618149316045
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011110110111010011111110;
 b = 32'b00111110110001110100111111001111;
 correct = 32'b00111110110000111100011001010110;
 #400 //0.9822539148219761 * 0.3892807614916026 = 0.38237255194000663
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001100011001101100011111;
 b = 32'b00111111011101110110101011000000;
 correct = 32'b00111111001010111010011010111010;
 #400 //0.6937731938729998 * 0.9664725981317817 = 0.6705127811966224
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110010010111101010111000;
 b = 32'b00111110001000001000111100100010;
 correct = 32'b00111101011111001011101010110010;
 #400 //0.3935143853294679 * 0.15679600905647795 = 0.06170148512597361
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110100011101101101010000011;
 b = 32'b00111110001111110011110010101001;
 correct = 32'b00111101010101010110110111000011;
 #400 //0.2790108631743913 * 0.1867548445646402 = 0.05210663038397954
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000100011110000000101000;
 b = 32'b00111111010111100001000001010110;
 correct = 32'b00111110111111010001001101100100;
 #400 //0.5698266172390777 * 0.8674367732156574 = 0.494288562150259
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010011110011001001000010;
 b = 32'b00111110101000111100100110011110;
 correct = 32'b00111110100001001001000000101110;
 #400 //0.8093606296061023 * 0.3198975890383505 = 0.2589125140735536
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110010001110000101011010100;
 b = 32'b00111111000111010110111000100101;
 correct = 32'b00111101111101001100111010001111;
 #400 //0.19437724046727578 * 0.6149619321060986 = 0.11953460335520766
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011001101000011111100011;
 b = 32'b00111111001010100001100101001100;
 correct = 32'b00111111000110010010110100000101;
 #400 //0.9005109655900614 * 0.6644485254870012 = 0.598343183271192
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110111000000100110010010110;
 b = 32'b00111111010000100011101110010011;
 correct = 32'b00111110101010100010111000111100;
 #400 //0.43808431620102917 * 0.7587215165724797 = 0.33238399677466257
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001100001101101001101110;
 b = 32'b00111111000101100100000001101000;
 correct = 32'b00111110110011111001100011110110;
 #400 //0.6908329933654739 * 0.5869202495589726 = 0.405463872869636
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000010101111010100001011;
 b = 32'b00111110111100110011100011101110;
 correct = 32'b00111110100001000000010110000000;
 #400 //0.5428015665389455 * 0.47504369935575563 = 0.25785446418476005
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101100110000101101100001010;
 b = 32'b00111110101100110100000000010010;
 correct = 32'b00111100110101010101101110010011;
 #400 //0.07439239541513332 * 0.35009819275441434 = 0.026044643189509952
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111000101010000101011001110;
 b = 32'b00111101100011100000101110000101;
 correct = 32'b00111101001001010110010101100110;
 #400 //0.5821961203229079 * 0.0693579059298367 = 0.040379903746072136
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010111101001110000010111;
 b = 32'b00111111010100011101010110110111;
 correct = 32'b00111111001101100111011101000110;
 #400 //0.8695692348979237 * 0.8196672687489424 = 0.7127574397568887
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110000011111111100010111;
 b = 32'b00111110001110110111011111001000;
 correct = 32'b00111101100011100001000000011011;
 #400 //0.37889931097410445 * 0.18307412108421217 = 0.06936665833599776
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110111100100011001011010000;
 b = 32'b00111111001101010100100100111000;
 correct = 32'b00111110101010111000001100110011;
 #400 //0.473043909995566 * 0.7081484919228349 = 0.33498533147664133
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011100101010010001101101;
 b = 32'b00111111011110010010000001000100;
 correct = 32'b00111111011011000010000010000011;
 #400 //0.9478214149812183 * 0.973148592691786 = 0.9223710761121099
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111101011101101010001100100100;
 b = 32'b00111101100001110111101011000101;
 correct = 32'b00111011100000101000011001001111;
 #400 //0.060214177986228634 * 0.06615213097765271 = 0.003983296188856689
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111001101110001101110010110;
 b = 32'b00111111000000111101100100011000;
 correct = 32'b00111110101111001001110011001001;
 #400 //0.715264651217978 * 0.5150313088723972 = 0.3683836895069539
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010001000000011000110101;
 b = 32'b00111111000000010100101000011001;
 correct = 32'b00111110110001011111111110111100;
 #400 //0.7657197181686372 * 0.5050368995403881 = 0.3867167123808283
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110010100001101010111110011;
 b = 32'b00111110101101001110100011110111;
 correct = 32'b00111101100100111001010001111010;
 #400 //0.20394114771545746 * 0.3533398866256868 = 0.0720605420120922
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110111000010001000101001;
 b = 32'b00111110101101100001101011100100;
 correct = 32'b00111110000111001001011101101000;
 #400 //0.42994810970967934 * 0.35567390905400076 = 0.15292132487082002
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011010110100010110010100;
 b = 32'b00111111010111110111100111000001;
 correct = 32'b00111111010011010110000110000001;
 #400 //0.9190304078264891 * 0.8729515969365622 = 0.8022690621453937
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110101010011111001110000101;
 b = 32'b00111111010011001011110100110001;
 correct = 32'b00111110100001111110101110100111;
 #400 //0.33193602331115624 * 0.7997618532645832 = 0.2654697691686062
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111011110101110101011001110;
 b = 32'b00111111011110010001011101100110;
 correct = 32'b00111111011101000010010101010010;
 #400 //0.9801453323235508 * 0.973013295663074 = 0.9536944400329171
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010011100000100000100101;
 b = 32'b00111110101000000100111010100010;
 correct = 32'b00111110100000010000010001100000;
 #400 //0.80481179416883 * 0.3130999247037991 = 0.2519865121549901
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110101001100110100100101011;
 b = 32'b00111101111001000001010111100010;
 correct = 32'b00111101000101000100001111100011;
 #400 //0.3250211042793112 * 0.11136986159487239 = 0.03619755539899947
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110001010111110110010101011;
 b = 32'b00111111000001110110000010111111;
 correct = 32'b00111101101101011101010110001111;
 #400 //0.16789500475982866 * 0.528820002981106 = 0.0887862369176054
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111110110010111001101110111111;
 b = 32'b00111110100000001100010011011100;
 correct = 32'b00111101110011001101010011100011;
 #400 //0.3976726092393811 * 0.25150192592630294 = 0.10001542711184243
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end

 a = 32'b00111111010101110111000111111011;
 b = 32'b00111111000011000000111010000000;
 correct = 32'b00111110111010111011110100010011;
 #400 //0.841582933773089 * 0.5470962723513849 = 0.4604268859417994
 if ((correct - out > 2) && (out - correct > 2)) begin
 $display ("A     : %b B      : %b", a, b);
 $display ("Output: %b Correct: %b", out, correct); end
 $finish;
 // stop the simulation
 end

endmodule
