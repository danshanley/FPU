//-----------------------------------------------------------
// File: fpu_tb.v
// FPU Test Bench
//-----------------------------------------------------------
`timescale 1 ns/100 ps
module fpu_tb ();
 //----------------------------------------------------------
 // inputs to the DUT are reg type
 reg clock;
 reg [31:0] a, b;
 reg [1:0] op;
 reg [31:0] correct;
 //----------------------------------------------------------
 // outputs from the DUT are wire type
 wire [31:0] out;
 wire [49:0] pro;
 //----------------------------------------------------------
 // instantiate the Device Under Test (DUT)
 // using named instantiation
 fpu U1 (
          .clk(clock),
          .A(a),
          .B(b),
          .opcode(op),
          .outp(out)
        );
 //----------------------------------------------------------
 // create a 10Mhz clock
 always
 #100 clock = ~clock; // every 100 nanoseconds invert
 //----------------------------------------------------------
 // initial blocks are sequential and start at time 0
 initial
 begin
 $dumpfile("fpu_tb.vcd");
 $dumpvars(0,clock, a, b, op, out);
 clock = 0;op = 2'b01;
a = 32'b00111111001000100000011101101100;
b = 32'b00111110111010110111001010010111;
correct = 32'b00111110001100010011100010000001;
#400 //0.632925725975876 * 0.45985861330843436 = 0.17306711266744168
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000011011010000011000001;
b = 32'b00111110110111010011010000011101;
correct = 32'b00111101111110000011010110010010;
#400 //0.5532341406472623 * 0.4320382122911741 = 0.12119592835608817
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010000000011010101110100;
b = 32'b00111111001000011101111010011001;
correct = 32'b00111101111100101011011011010111;
#400 //0.7508156110895009 * 0.632302808425902 = 0.11851280266359887
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110111001010101011010111000;
b = 32'b00111110111011111000111110111010;
correct = 32'b10111100101000111001000000010101;
#400 //0.4479272483332768 * 0.4678934133281276 = -0.01996616499485082
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110010000001010110011000001;
b = 32'b00111111011001000100010100010011;
correct = 32'b10111111001101000001100111100011;
#400 //0.18815900418327158 * 0.8916789780943901 = -0.7035199739111185
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010000101000111110011100;
b = 32'b00111111010011011000011101011010;
correct = 32'b10111101001011110111101111100101;
#400 //0.7600037989237857 * 0.802846561597781 = -0.04284276267399534
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101011000011111000110011;
b = 32'b00111111011001111100110111011110;
correct = 32'b10111111000100011010111011000100;
#400 //0.3364120339027663 * 0.9054850112100754 = -0.5690729773073091
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101010111110101100011011;
b = 32'b00111110111000001110110010101001;
correct = 32'b10111101110101000000011000110110;
#400 //0.33577810090755944 * 0.43930557177209173 = -0.10352747086453229
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101111000010111001001001010;
b = 32'b00111111000001011100101110011110;
correct = 32'b10111110110100110011101010101010;
#400 //0.11008126992720701 * 0.5226382184408391 = -0.4125569485136321
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100001101000011010010000;
b = 32'b00111111011010000010010011001100;
correct = 32'b10111111001001001110000110000100;
#400 //0.26274538909186596 * 0.9068114946553414 = -0.6440661055634754
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001111010010001001111111;
b = 32'b00111111011001000111111011000111;
correct = 32'b10111110000111010111000100011110;
#400 //0.7388076164170791 * 0.8925594394637497 = -0.15375182304667057
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001011110000011100001001;
b = 32'b00111101110010100110111010001111;
correct = 32'b00111111000101011011100100111000;
#400 //0.6837011201108391 * 0.09884368518403264 = 0.5848574349268064
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101111110101000100011110000;
b = 32'b00111110110001001111010111100011;
correct = 32'b10111110100001100101001110100111;
#400 //0.12233149842213753 * 0.38468847399947026 = -0.26235697557733273
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101101010110011101000001100;
b = 32'b00111110110110111101111000101000;
correct = 32'b10111110101100010000111110100101;
#400 //0.08360681296105466 * 0.42942930627222475 = -0.3458224933111701
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110110110010010101100000;
b = 32'b00111110011000000000110010101111;
correct = 32'b00111110010101100011111000010010;
#400 //0.4280195356856642 * 0.21879838492456782 = 0.20922115076109637
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110111110000101001010010011;
b = 32'b00111111010011010100110001110101;
correct = 32'b10111110101000100100011001011000;
#400 //0.48500498600502273 * 0.8019479153698578 = -0.31694292936483504
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110010100001100111000001110;
b = 32'b00111111010100011011001111110110;
correct = 32'b10111111000111011000000001110010;
#400 //0.2039110311337483 * 0.819152219196945 = -0.6152411880631967
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110001110010100110010011;
b = 32'b00111111011000001111010011110100;
correct = 32'b10111110111110101100000001010100;
#400 //0.388989075046525 * 0.8787376726091192 = -0.48974859756259415
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110001101100001110000100110;
b = 32'b00111110000101100001011010011001;
correct = 32'b00111101000000000001011000110011;
#400 //0.17784174758263016 * 0.1465705749283791 = 0.031271172654251056
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100100111100111001110101;
b = 32'b00111101100101011000000110011100;
correct = 32'b00111110010111001101110000011100;
#400 //0.2886845210411898 * 0.07300111411122256 = 0.21568340692996724
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001011011001011110010000;
b = 32'b00111111001110000010001000011110;
correct = 32'b10111101001010001010100011100111;
#400 //0.6780938879735791 * 0.7192705898584137 = -0.04117670188483469
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010100110000011000001100;
b = 32'b00111110101100001011100010001101;
correct = 32'b00111110111101010101001110001100;
#400 //0.82431104237697 * 0.3451579995058549 = 0.47915304287111504
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100011001000000001001110;
b = 32'b00111110001001011010000010010111;
correct = 32'b00111101111001101100000000001100;
#400 //0.27441639144509555 * 0.16174540720364017 = 0.11267098424145539
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101101111100100000111011110;
b = 32'b00111111010011111111100101110000;
correct = 32'b10111111001110000011000100110100;
#400 //0.09289906754486232 * 0.8123998479920311 = -0.7195007804471688
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101111111010101101010011100;
b = 32'b00111111000101000000011000101111;
correct = 32'b10111110111010001011010110110111;
#400 //0.12370798309755571 * 0.5782193688588704 = -0.45451138576131467
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011011100001001111100000;
b = 32'b00111111001000000100000001010101;
correct = 32'b00111110100110111010011100010110;
#400 //0.9299907861259514 * 0.6259816345097992 = 0.3040091516161523
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101000001111101111111100000;
b = 32'b00111110100011011101111001100100;
correct = 32'b10111110011110011100010011010001;
#400 //0.03317248927006311 * 0.27708734057239515 = -0.24391485130233204
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101100100100101010001110;
b = 32'b00111110010010111110001001110010;
correct = 32'b00111110000110001011001010101011;
#400 //0.34822507086721777 * 0.1991060031906582 = 0.14911906767655958
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110111101101001011110110101;
b = 32'b00111111011011110101000101101101;
correct = 32'b10111110111010000000101100100101;
#400 //0.48162618695977955 * 0.9348362176156173 = -0.45321003065583776
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010110011001110101100010;
b = 32'b00111111000000011001001000000100;
correct = 32'b00111110101100000001011010111100;
#400 //0.8500577494493873 * 0.5061342886663501 = 0.34392346078303715
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110000111011010010101111111;
b = 32'b00111110110010111100110011110000;
correct = 32'b10111110011110011111010001100000;
#400 //0.153951635758371 * 0.3980479203535714 = -0.24409628459520039
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101010100001000110011100;
b = 32'b00111110010010011110000111100001;
correct = 32'b00111110000010100100000101010111;
#400 //0.33216560450624655 * 0.197150727982355 = 0.13501487652389155
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011110011000010110010010;
b = 32'b00111110111010010100100110011100;
correct = 32'b00111111000001001110000011000100;
#400 //0.9746943911441196 * 0.4556397311789582 = 0.5190546599651614
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010110101111100100001100;
b = 32'b00111111001000100110011100000000;
correct = 32'b00111110011000100100100000110001;
#400 //0.8553626830836216 * 0.634384175784475 = 0.2209785072991466
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000000111100011011001110;
b = 32'b00111111010101001100010111010100;
correct = 32'b10111110101000011111111000001100;
#400 //0.5147522478131229 * 0.8311436078729016 = -0.31639136005977875
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010001110110101001001111;
b = 32'b00111111011101110100011111011000;
correct = 32'b10111110001111110111011000100101;
#400 //0.7789658992538196 * 0.9659400165986657 = -0.18697411734484604
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010111101011100011010000;
b = 32'b00111111001001110011000010100011;
correct = 32'b00111110010111100010000010110110;
#400 //0.8700075250025203 * 0.6530858680770426 = 0.2169216569254777
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110111110011101110001011000;
b = 32'b00111111011111001100100111001101;
correct = 32'b10111110111111111011011101000010;
#400 //0.48800921589352975 * 0.9874542463312178 = -0.49944503043768806
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110110011010001110111110;
b = 32'b00111111001101111010110101010111;
correct = 32'b10111110100101011011011011101111;
#400 //0.42507736805685414 * 0.7174886773870144 = -0.29241130933016024
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011110001110011111111010;
b = 32'b00111101001100001010111110101001;
correct = 32'b00111111011011011101110100000000;
#400 //0.9722896919753771 * 0.04313627404748699 = 0.9291534179278901
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010010111100110011000111;
b = 32'b00111110100011111101011011101000;
correct = 32'b00111111000000111110000101010011;
#400 //0.7960934070581507 * 0.2809364856724266 = 0.5151569213857241
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001101011110001011111000;
b = 32'b00111111001101010011111000100100;
correct = 32'b00111011001001001101001111100001;
#400 //0.7104945254228882 * 0.7079794551506509 = 0.0025150702722372964
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100011110110010100101111;
b = 32'b00111111001110010111010001100110;
correct = 32'b10111110111000111000001110011100;
#400 //0.28006885413976956 * 0.724432320804853 = -0.4443634666650834
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010000101010001110001110;
b = 32'b00111111010000000111010000110001;
correct = 32'b00111100000010111101011100001110;
#400 //0.7603081222050291 * 0.7517729623437436 = 0.008535159861285502
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001100000011110000111001;
b = 32'b00111111000000010011111101110011;
correct = 32'b00111110001110111111001100011001;
#400 //0.688418942839271 * 0.504874416778359 = 0.18354452606091198
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110011011110101001011100111;
b = 32'b00111111000001110011011100011011;
correct = 32'b10111110100101101100010011000010;
#400 //0.23371468594515743 * 0.5281845712278459 = -0.29446988528268847
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010100111110100100000001;
b = 32'b00111110111101110001000011100110;
correct = 32'b00111110101100001100000100011100;
#400 //0.8277741033216073 * 0.4825508025270169 = 0.3452233007945904
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011001111010011011111001;
b = 32'b00111110010011001111011010101100;
correct = 32'b00111111001101000110100101001110;
#400 //0.9048915580522362 * 0.20015973503047768 = 0.7047318230217585
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110011111000111101100101;
b = 32'b00111110100111111100001011011110;
correct = 32'b00111101101111110011001000011101;
#400 //0.4053908825736595 * 0.3120335823430763 = 0.0933573002305832
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000010101110010000101111;
b = 32'b00111110101110000010000100110011;
correct = 32'b00111110001110110100111001010110;
#400 //0.5425443121255309 * 0.3596282954996486 = 0.1829160166258823
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110001101110000001110101;
b = 32'b00111111000110110000100000000011;
correct = 32'b10111110010111100101111100100001;
#400 //0.3884312297359668 * 0.6055909901580832 = -0.21715976042211638
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001101110110101010011110;
b = 32'b00111111001110011000101000111011;
correct = 32'b10111100000001111110011100111111;
#400 //0.7164706138951633 * 0.7247654936919932 = -0.008294879796829857
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010010010010101010010001;
b = 32'b00111111000010100111010011010101;
correct = 32'b00111110011110101101011011110001;
#400 //0.7858057570332081 * 0.540845195904802 = 0.24496056112840614
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101001000100001001110001110;
b = 32'b00111111010111010101010001010001;
correct = 32'b10111111010100110011001100011000;
#400 //0.03956942847580003 * 0.8645678089014927 = -0.8249983804256926
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010001010111011011101111;
b = 32'b00111111010000110001101010000000;
correct = 32'b00111100000101110001101111010101;
#400 //0.7713460505568208 * 0.7621231065729395 = 0.009222943983881349
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110111010110110010100110001;
b = 32'b00111110001010011000110000110001;
correct = 32'b00111110100101101001111100011000;
#400 //0.45975639059093754 * 0.16557385174443373 = 0.2941825388465038
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001001011000000101010001;
b = 32'b00111110110010111000110111111110;
correct = 32'b00111110011111101110100101001000;
#400 //0.6465044553929735 * 0.3975676800767024 = 0.24893677531627112
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010011110110010101011000;
b = 32'b00111111010011001011100011000000;
correct = 32'b00111100001010110010011000000010;
#400 //0.8101401455705267 * 0.7996940723799847 = 0.010446073190542027
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001000101000010001011111;
b = 32'b00111110000000010001100001101110;
correct = 32'b00111111000000100011111001000011;
#400 //0.6348322929740232 * 0.1260697557838074 = 0.5087625371902158
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000000100010101000001010;
b = 32'b00111110011011111100011110011010;
correct = 32'b00111110100011000111000001000111;
#400 //0.5084539574210768 * 0.23415985335482914 = 0.27429410406624766
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100000001101110110010110;
b = 32'b00111101111100110100101110011110;
correct = 32'b00111110000010000001010101011100;
#400 //0.25169055414637065 * 0.11879657250089826 = 0.1328939816454724
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011101111001100100111010;
b = 32'b00111101101110000110000011111110;
correct = 32'b00111111011000001000110100011010;
#400 //0.9671817904529433 * 0.09002874771992964 = 0.8771530427330136
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011111110000000010101010;
b = 32'b00111110101001111111011001110011;
correct = 32'b00111111001010110000010101110000;
#400 //0.9961038623424072 * 0.32805211995983297 = 0.6680517423825743
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101110001111011011101111;
b = 32'b00111111010010011111011100001100;
correct = 32'b10111110110110101111011100101001;
#400 //0.36125894400726266 * 0.7889258631655689 = -0.42766691915830624
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110000010100010000001000011;
b = 32'b00111110000110110101001001111010;
correct = 32'b10111100100010011001000110110101;
#400 //0.13488869744624987 * 0.15168180936918252 = -0.016793111922932646
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000101110011111011100001;
b = 32'b00111111000110110010101100110101;
correct = 32'b10111100011110110001010011100100;
#400 //0.5908032222011934 * 0.6061280274218018 = -0.015324805220608417
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000000010010010010101111;
b = 32'b00111110100000001111110111000100;
correct = 32'b00111110100000010100101110011010;
#400 //0.5044660056179193 * 0.2519360905043754 = 0.25252991511354395
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011011100010001010101001;
b = 32'b00111111010011001011101010110000;
correct = 32'b00111110000001011001111111100111;
#400 //0.9302163935973401 * 0.7997235971704587 = 0.13049279642688139
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000101010100011101000110;
b = 32'b00111110111101011010111110010111;
correct = 32'b00111101110100110111101111010010;
#400 //0.5831187878793451 * 0.47985527503171777 = 0.10326351284762736
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011000010110100100001111;
b = 32'b00111110100000010000111100110001;
correct = 32'b00111111001000001110000101110110;
#400 //0.8805092971163266 * 0.2520690388500457 = 0.6284402582662809
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101000111011100110011111;
b = 32'b00111111001001001101001000011101;
correct = 32'b10111110101001011110101010011011;
#400 //0.3197755640376737 * 0.6438310811101824 = -0.3240555170725087
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001011010001101011010110;
b = 32'b00111111000100011000011011001010;
correct = 32'b00111101110111001010000001011111;
#400 //0.6761907485129671 * 0.5684629898906884 = 0.10772775862227868
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110111100101100001000101111;
b = 32'b00111111011010010101110010110011;
correct = 32'b10111110110111111111011100110110;
#400 //0.47413776088636117 * 0.9115707156176941 = -0.4374329547313329
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101110111100100010100111010;
b = 32'b00111111001011111011110001000111;
correct = 32'b10111111000100111111001110011111;
#400 //0.1085304752807923 * 0.6864666078443608 = -0.5779361325635685
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101000010010010111000010;
b = 32'b00111110011000111011100011000011;
correct = 32'b00111101101111010010010110000011;
#400 //0.3147412005635444 * 0.22238449910997393 = 0.09235670145357044
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101100110110010011001101;
b = 32'b00111110010110000001010111111111;
correct = 32'b00111110000011101011001110011010;
#400 //0.35037842254025275 * 0.21102141552291842 = 0.13935700701733433
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101011100100111100111100111;
b = 32'b00111111001000001110100100011100;
correct = 32'b10111111000100011100000101111110;
#400 //0.0591982874528072 * 0.628556991328566 = -0.5693587038757588
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101110111100111010110110;
b = 32'b00111110011111111011000011110100;
correct = 32'b00111101111011111101100011110000;
#400 //0.36681146039076107 * 0.24969846690718567 = 0.1171129934835754
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100101100101010000000100;
b = 32'b00111111010110001001110101100110;
correct = 32'b10111111000011010111001101100100;
#400 //0.2936097237596609 * 0.8461517094403658 = -0.5525419856807049
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111100100010110010011100110100;
b = 32'b00111111010011110010111011100011;
correct = 32'b10111111010010101101010110101001;
#400 //0.016986466395788713 * 0.8093091891653883 = -0.7923227227695996
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110000110100111110100101100;
b = 32'b00111111001111100100011100110111;
correct = 32'b10111111000101111010011111101100;
#400 //0.15086811501302044 * 0.7432741714323823 = -0.5924060564193618
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110000101100111010000100100;
b = 32'b00111111001011001000110110101110;
correct = 32'b10111111000001101111000010100101;
#400 //0.14692741220640637 * 0.6740368446002933 = -0.527109432393887
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111011111010111110010000111001;
b = 32'b00111111011010110110111111011001;
correct = 32'b10111111011010011001100000010001;
#400 //0.007198836910069284 * 0.9196754366747368 = -0.9124765997646676
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001100100000101111011001;
b = 32'b00111111011011100111010111010111;
correct = 32'b10111110011100011010011111111011;
#400 //0.695493262895544 * 0.9314856138001179 = -0.23599235090457382
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110001001110000000011000;
b = 32'b00111110000100111010001101011111;
correct = 32'b00111110011101100001110011010001;
#400 //0.38452219511637753 * 0.14417789640315015 = 0.24034429871322738
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100101001000111110110100;
b = 32'b00111111001111100100110100011001;
correct = 32'b10111110111010000000101001111110;
#400 //0.29015886404202595 * 0.7433639270110168 = -0.4532050629689909
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100100011011001101001000;
b = 32'b00111111000001100111110010011110;
correct = 32'b10111110011101101000101111100110;
#400 //0.28457093916041976 * 0.5253389834298386 = -0.2407680442694189
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100001010001001111010110;
b = 32'b00111110011010000111010100111110;
correct = 32'b00111101000001101100100110110111;
#400 //0.25991695986240615 * 0.22700974668274831 = 0.032907213179657835
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111101010011111011001111100110;
b = 32'b00111110111110011100101000100101;
correct = 32'b10111110110111111101001110101000;
#400 //0.05070867414506197 * 0.4878703680148958 = -0.43716169386983383
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110101110100111110010101111;
b = 32'b00111100111010111111101010010101;
correct = 32'b00111110101010111011110100000110;
#400 //0.36423251746596996 * 0.028806009658597587 = 0.3354265078073724
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110101101011010011011100;
b = 32'b00111111011110000010011111000100;
correct = 32'b10111111000011001100110101010101;
#400 //0.41934860989013734 * 0.9693567561924049 = -0.5500081463022676
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010000111101101111010010;
b = 32'b00111111011010010011101001000010;
correct = 32'b10111110000101010111100111000010;
#400 //0.7650729388437663 * 0.9110452197364639 = -0.14597228089269765
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111010101010001100010000000;
b = 32'b00111101100101111111010100101010;
correct = 32'b00111111010000100001100111011010;
#400 //0.8324050748358335 * 0.07419808526283356 = 0.7582069895729999
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110100100000000010100101000;
b = 32'b00111110000010101101001001010111;
correct = 32'b00111110000101010011011111111001;
#400 //0.2812893303317834 * 0.13556800579839456 = 0.14572132453338882
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110010111001111011011111011;
b = 32'b00111111010000100111101011011000;
correct = 32'b10111111000010110011110100011001;
#400 //0.21578590791836094 * 0.7596869353928337 = -0.5439010274744728
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000011010011110101111010;
b = 32'b00111110010000110010001111100001;
correct = 32'b00111110101110001110100100000011;
#400 //0.5517192941585503 * 0.19056655891964636 = 0.3611527352389039
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111001110100100111000011101;
b = 32'b00111111000110111111001111000011;
correct = 32'b00111101111100101101001011001100;
#400 //0.727754407219723 * 0.6091882793076714 = 0.11856612791205157
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111011011110100100010110001;
b = 32'b00111110101001101011100111101000;
correct = 32'b00111111000110111110101110111101;
#400 //0.9347029435607085 * 0.32563710000010415 = 0.6090658435606043
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111111000010111011000111110011;
b = 32'b00111111000110100111000001010011;
correct = 32'b10111101011010111110011000000101;
#400 //0.5456840192153833 * 0.603276431032947 = -0.05759241181756369
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
a = 32'b00111110110101111011100100101001;
b = 32'b00111110001100010010000010101011;
correct = 32'b00111110011111100101000110100111;
#400 //0.4213345348845866 * 0.17297618596567366 = 0.24835834891891295
if (correct[31:11] != out[31:11]) begin
$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
$display ("Correct: %b %b %b",correct[31], correct[30:23], correct[22:0]); end
$display ("Done.");
$finish;
 // stop the simulation
 end

endmodule